package datatypes;
import FixedPoint::*;
typedef FixedPoint#(10,6) DataType;
typedef UInt#(16) ImgWidth;
typedef FixedPoint#(2,14) CoeffType;
typedef UInt#(9) Width;
typedef Bit#(16) Tin;
typedef Int#(16) Tin2;

endpackage
